module control
#(
    // Parameters.

)
(
    // Outputs.

    // Inputs.

) ;

    //==========================================================================
    // LOCAL PARAMETERS.
    //==========================================================================


    //==========================================================================
    // INTERNAL SIGNALS.
    //==========================================================================

    //==========================================================================
    // ALGORITHM.
    //==========================================================================

endmodule